`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    12:19:21 04/15/2016 
// Design Name: 
// Module Name:    CPU_SameDickNewBush 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module CPU_SameDickNewBush(
    );
	 
	 CPU_Datapath JebBush ();
	 CPU_Control DickChaney();


endmodule
